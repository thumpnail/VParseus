module ebnf_ast

