module ebnf
fn parser() {

}