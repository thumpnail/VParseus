module ebnf
fn lexer() {

}