module ebnf

fn (mut ctx VParseusContext)build_parser(node SyntaxNode) string {
	code := ""
	return code
}
