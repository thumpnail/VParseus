module ebnf

fn (mut ctx VParseusContext)build_ast_structure(node SyntaxNode) string {
	code := ""
	return code
}
