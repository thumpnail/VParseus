module ebnf

pub fn (mut ctx VParseusContext) finalize(ebnf_path string, token_path string) {}
