module scretches
