module scretches

fn preprocessor() []string {
// start := { stat };
//stat := data_decl
//    | assign
//    | decl;
//data_decl := 'data' { expr_list } '{' decl '}';
//assign := identifier [ ':' type ] := expr;
//decl := identifier [ ':' type ];
//expr := expr | expr '+' expr | expr '*' expr | number;
//expr_list := expr { ',' expr };
//identifier := '[a-zA-Z_0-9]';
//number := ['-'] '[0-9]+';
}
